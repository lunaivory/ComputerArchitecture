//TODO
module Hazard_Detection_Unit(
  input       [31:0]  inst_i,
  input       [4:0]   IDEX_RT_addr_i,
  input               IDEX_MemRead_i,
  output reg  [31:0]  PC_o,
  output reg          IF_ID_o,
  output reg          flush_o
);

endmodule