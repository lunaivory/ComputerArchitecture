//TODO
module Data_Memory(
  input             clk_i,
  input      [31:0] addr_i,
  input      [31:0] write_data_i,
  input             MemRead_i,
  input             MemWrite_i,
  output reg [31:0] data_o
);

endmodule