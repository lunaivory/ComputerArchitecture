//TODO
module Equal(
  input [31:0] data1_i,
  input [31:0] data2_i,
  output reg   data_o
);
endmodule