//TODO
module ForwardMUX(
  input      [31:0] data0_i,
  input      [31:0] data1_i,
  input      [31:0] data2_i,
  input      [1:0]  select_i,
  output reg [31:0] data_o
);

endmodule