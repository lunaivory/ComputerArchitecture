//TODO
module Shift_Left2_Concat(
  input       [25:0]  inst_i,
  input       [3:0]   addedPC_i,
  output reg  [31:0]  jumpAddr_o
);

endmodule