//TODO
module Shift_Left2(
  input      [31:0] data_i,
  output reg [31:0] data_o
);

endmodule