//NOT MODIFIED
module Signed_Extend(
  input   [15:0]  data_i,
  output  [31:0]  data_o
);
assign data_o = data_i;

endmodule