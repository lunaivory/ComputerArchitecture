//TODO
module Flush_MUX(
  input      [1:0]  WB_i,
  input      [2:0]  EX_i,
  input      [1:0]  MEM_i,
  input             flush_i,
  output reg [1:0]   WB_o,
  output reg [2:0]  EX_o,
  output reg [1:0]  MEM_o 
);

endmodule